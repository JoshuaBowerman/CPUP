`timescale 1ns / 1ps

module memory_controller(
output 			ras,
output 			cas,
output			we,
output			oe,
output [12:0]	dram_addr,
inout  [15:0]	dram_dq,
inout  [15:0]	bus,
input  [15:0]	address_space,
input  [2:0]	mem_control_bus,
input				clock

);





endmodule 